module Segmentos(input logic bcd, output logic [6:0] seg,seg2);
//acá hay que hacerlo para 6 bits, es decir hasta el 63
  always_comb begin 
    case (bcd)
		0: {seg, seg2} = {7'b0000001, 7'b0000000}; // numero 0
		1: {seg, seg2} = {7'b1001111, 7'b0000000}; // numero 1
		2: {seg, seg2} = {7'b0010010, 7'b0000000}; // numero 2
		3: {seg, seg2} = {7'b0000110, 7'b0000000}; // numero 3
		4: {seg, seg2} = {7'b1001100, 7'b0000000}; // num 4
		5: {seg, seg2} = {7'b0100100, 7'b0000000}; // num 5
		6: {seg, seg2} = {7'b0100000, 7'b0000000}; // num 6
		7: {seg, seg2} = {7'b0001111, 7'b0000000}; // num 7
		8: {seg, seg2} = {7'b0000000, 7'b0000000}; // num 8
		9: {seg, seg2} = {7'b0000100, 7'b0000000}; // num 9
		10: {seg, seg2} = {7'b0001000, 7'b0000000}; // A hex 10
		11: {seg, seg2} = {7'b1100000, 7'b0000000}; // B hex 11
		12: {seg, seg2} = {7'b0110001, 7'b0000000}; // C    12
		13: {seg, seg2} = {7'b1000010, 7'b0000000}; // D    13
		14: {seg, seg2} = {7'b0110000, 7'b0000000}; // E    14
		15: {seg, seg2} = {7'b0111000, 7'b0000000}; // F    15
		16: {seg, seg2} = {7'b0000001, 7'b1001111}; // 16
		17: {seg, seg2} = {7'b1001111, 7'b1001111}; // 17
		18: {seg, seg2} = {7'b0010010, 7'b1001111}; // 18
		19: {seg, seg2} = {7'b0000110, 7'b1001111}; // 19
		20: {seg, seg2} = {7'b1001100, 7'b1001111}; // 20
		21: {seg, seg2} = {7'b0100100, 7'b1001111}; // 21
		22: {seg, seg2} = {7'b0100000, 7'b1001111}; // 22
		23: {seg, seg2} = {7'b0001111, 7'b1001111}; // 23
		24: {seg, seg2} = {7'b0000000, 7'b1001111}; // 24
		25: {seg, seg2} = {7'b0000100, 7'b1001111}; // 25
		26: {seg, seg2} = {7'b0001000, 7'b1001111}; // 26
		27: {seg, seg2} = {7'b1100000, 7'b1001111}; // 27
		28: {seg, seg2} = {7'b0110001, 7'b1001111}; // 28
		29: {seg, seg2} = {7'b1000010, 7'b1001111}; // 29
		30: {seg, seg2} = {7'b0110000, 7'b1001111}; // 30
		31: {seg, seg2} = {7'b0111000, 7'b1001111}; // 31
		32: {seg, seg2} = {7'b0000001, 7'b0010010}; // 32
		33: {seg, seg2} = {7'b1001111, 7'b0010010}; // 33
		34: {seg, seg2} = {7'b0010010, 7'b0010010}; // 34
		35: {seg, seg2} = {7'b0000110, 7'b0010010}; // 35
		36: {seg, seg2} = {7'b1001100, 7'b0010010}; // 36
		37: {seg, seg2} = {7'b0100100, 7'b0010010}; // 37
		38: {seg, seg2} = {7'b0100000, 7'b0010010}; // 38
		39: {seg, seg2} = {7'b0001111, 7'b0010010}; // 39
		40: {seg, seg2} = {7'b0000000, 7'b0010010}; // 40
		41: {seg, seg2} = {7'b0000100, 7'b0010010}; // 41
		42: {seg, seg2} = {7'b0001000, 7'b0010010}; // 42
		43: {seg, seg2} = {7'b1100000, 7'b0010010}; // 43
		44: {seg, seg2} = {7'b0110001, 7'b0010010}; // 44
		45: {seg, seg2} = {7'b1000010, 7'b0010010}; // 45
		46: {seg, seg2} = {7'b0110000, 7'b0010010}; // 46
		47: {seg, seg2} = {7'b0111000, 7'b0010010}; // 47
		48: {seg, seg2} = {7'b0000001, 7'b0000110}; // 48
		49: {seg, seg2} = {7'b1001111, 7'b0000110}; // 49
		50: {seg, seg2} = {7'b0010010, 7'b0000110}; // 50
		51: {seg, seg2} = {7'b0000110, 7'b0000110}; // 51
		52: {seg, seg2} = {7'b1001100, 7'b0000110}; // 52
		53: {seg, seg2} = {7'b0100100, 7'b0000110}; // 53
		54: {seg, seg2} = {7'b0100000, 7'b0000110}; // 54
		55: {seg, seg2} = {7'b0001111, 7'b0000110}; // 55
		56: {seg, seg2} = {7'b0000000, 7'b0000110}; // 56
		57: {seg, seg2} = {7'b0000100, 7'b0000110}; // 57
		58: {seg, seg2} = {7'b0001000, 7'b0000110}; // 58
		59: {seg, seg2} = {7'b1100000, 7'b0000110}; // 59
		60: {seg, seg2} = {7'b0110001, 7'b0000110}; // 60
		61: {seg, seg2} = {7'b1000010, 7'b0000110}; // 61
		62: {seg, seg2} = {7'b0110000, 7'b0000110}; // 62
		63: {seg, seg2} = {7'b0111000, 7'b0000110}; // 63
			default: seg = 7'b1111111;
		endcase
	end
endmodule