module interfaz_tb();
endmodule;